module full_adder_no_tb();

	reg a,b,cin;
	wire sum,cout;

	full_adder_no FA1(a,b,cin,sum,cout);

	initial
	begin

	$monitor("Time=%t a=%b b=%b cin=%b sum=%b cout=%b",$time,a,b,cin,sum,cout);

	end
	initial
	begin

	 #0; {a,b,cin}=3'd0;
	#10; {a,b,cin}=3'd1;
	#10; {a,b,cin}=3'd2;
	#10; {a,b,cin}=3'd3;
	#10; {a,b,cin}=3'd4;
	#10; {a,b,cin}=3'd5;
	#10; {a,b,cin}=3'd6;
	#10; {a,b,cin}=3'd7;
	#10;
	$finish;

	end
endmodule

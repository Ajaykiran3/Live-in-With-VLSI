module full_subtractor_na(a,b,bin,diff,bout);

	input a,b,bin;
	output 	diff,bout;
	wire [6:0]w;

	nand NA1(w[0],a,b);
	nand NA2(w[1],a,w[0]);
	nand NA3(w[2],b,w[0]);
	nand NA4(w[3],w[1],w[2]);
	nand NA5(w[4],w[3],bin);
	nand NA6(w[5],w[3],w[4]);
	nand NA7(w[6],bin,w[4]);
	nand NA8(diff,w[5],w[6]);
	nand NA9(bout,w[2],w[6]);
endmodule
	

module decoder_2_4(
	input e,
	input [1:0]i,
	output reg [3:0]y);
	always@(i,e)
	begin
	if (e) begin
	case(i)
	2'd0:y=4'd1;
	2'd1:y=4'd2;
	2'd2:y=4'd4;
	2'd3:y=4'd8;
	default:y=2'bxx;
	endcase
	end
	else y=2'bxx;
	end
endmodule
module pri_enc_4_2(
	input [3:0]i,
	output reg [1:0]y);
	always@(i)
	begin
	casex(i)
	4'b0001:y=2'd0;
	4'b001x:y=2'd1;
	4'b01xx:y=2'd2;
	4'b1xxx:y=2'd3;
	default:y=2'bxx;
	endcase
	end
endmodule
